-- -*- vhdl -*-

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------
entity Division10 is
  port (
    rst         : in std_logic;
    clk         : in std_logic;
    clkDiv10    : out std_logic
    );
end Division10;

architecture RTL of Division10 is
  signal clk_inv  : std_logic;
  signal q_jk     : std_logic_vector(3 downto 0);
  signal in_jk    : std_logic_vector(3 downto 0);

  component JKFF is
    port(
      ACLR   : in std_logic;
      J	   : in std_logic;
      K      : in std_logic;
      CLK    : in std_logic;
      Q      : out std_logic
      );
  end component;

begin
  clkDiv10    <= q_jk(3);
  clk_inv     <= NOT clk;
  in_jk(0)    <= '1';
  in_jk(1)    <= q_jk(0) AND (NOT q_jk(3));
  in_jk(2)    <= q_jk(0) AND q_jk(1);
  in_jk(3)    <= (q_jk(0) AND q_jk(1) AND q_jk(2)) OR (q_jk(0) AND q_jk(3));

  gen_jkff : for i in 0 to 3 generate
    u_JK : JKFF
      port map(ACLR=>rst, J=>in_jk(i), K=>in_jk(i), CLK=>clk_inv, Q=>q_jk(i));
  end generate;
end RTL;
